module network_engine
(
    input logic CLK,
    input logic RST
);
    initial begin 
        $display("Hello World");
        $finish;
    end

endmodule 