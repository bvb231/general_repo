module mac_phy (
    input logic CLK
);

endmodule
