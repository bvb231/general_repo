module network_decoder
(
    input logic CLK, 
    input logic RST
);

endmodule